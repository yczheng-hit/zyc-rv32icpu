module bubble(
    input logic en
);
    
endmodule